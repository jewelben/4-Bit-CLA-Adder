* 5 Input AND gate
.subckt and5 OUT A B C D E 

*PUN
M0 5nand A vdd vdd CMOSP W={width_P} L={LAMBDA} +
AS={5*width_P*LAMBDA} PS={10*LAMBDA+2*width_P}
AD={5*width_P*LAMBDA} PD={10*LAMBDA+2*width_P}

M1 5nand B vdd vdd CMOSP W={width_P} L={LAMBDA} +
AS={5*width_P*LAMBDA} PS={10*LAMBDA+2*width_P}
AD={5*width_P*LAMBDA} PD={10*LAMBDA+2*width_P}

M2 5nand C vdd vdd CMOSP W={width_P} L={LAMBDA} +
AS={5*width_P*LAMBDA} PS={10*LAMBDA+2*width_P}
AD={5*width_P*LAMBDA} PD={10*LAMBDA+2*width_P}

M3 5nand D vdd vdd CMOSP W={width_P} L={LAMBDA} +
AS={5*width_P*LAMBDA} PS={10*LAMBDA+2*width_P}
AD={5*width_P*LAMBDA} PD={10*LAMBDA+2*width_P}

M4 5nand E vdd vdd CMOSP W={width_P} L={LAMBDA} +
AS={5*width_P*LAMBDA} PS={10*LAMBDA+2*width_P}
AD={5*width_P*LAMBDA} PD={10*LAMBDA+2*width_P}

*PDN
M5 5nand A node1 gnd CMOSN W={width_N} L={LAMBDA} +
AS={5*width_N*LAMBDA} PS={10*LAMBDA+2*width_N}
AD={5*width_N*LAMBDA} PD={10*LAMBDA+2*width_N}

M6 node1 B node2 gnd CMOSN W={width_N} L={LAMBDA} +
AS={5*width_N*LAMBDA} PS={10*LAMBDA+2*width_N}
AD={5*width_N*LAMBDA} PD={10*LAMBDA+2*width_N}

M7 node2 C node3 gnd CMOSN W={width_N} L={LAMBDA} +
AS={5*width_N*LAMBDA} PS={10*LAMBDA+2*width_N}
AD={5*width_N*LAMBDA} PD={10*LAMBDA+2*width_N}

M8 node3 D gnd node4 CMOSN W={width_N} L={LAMBDA} +
AS={5*width_N*LAMBDA} PS={10*LAMBDA+2*width_N}
AD={5*width_N*LAMBDA} PD={10*LAMBDA+2*width_N}

M9 node4 A gnd gnd CMOSN W={width_N} L={LAMBDA} +
AS={5*width_N*LAMBDA} PS={10*LAMBDA+2*width_N}
AD={5*width_N*LAMBDA} PD={10*LAMBDA+2*width_N}

*Inverter
M10 OUT 5nand VDD VDD CMOSP W={width_P} L={LAMBDA} +
AS={5*width_P*LAMBDA} PS={10*LAMBDA+2*width_P}
AD={5*width_P*LAMBDA} PD={10*LAMBDA+2*width_P}

M11 OUT 5nand GND Gnd CMOSN W={width_N} L={LAMBDA} +
AS={5*width_N*LAMBDA} PS={10*LAMBDA+2*width_N}
AD={5*width_N*LAMBDA} PD={10*LAMBDA+2*width_N}

.ends
