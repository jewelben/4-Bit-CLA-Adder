magic
tech scmos
timestamp 1638790149
<< metal1 >>
rect 243 665 359 670
rect 276 637 283 652
rect 262 632 283 637
rect -102 624 119 631
rect -103 616 165 621
rect 298 545 304 614
rect 262 540 304 545
rect 353 543 359 665
rect 938 559 946 567
rect -102 532 94 539
rect -103 524 165 529
rect 326 510 364 514
rect 326 509 331 510
rect 340 501 402 505
rect 340 500 345 501
rect 1142 464 1219 468
rect 1020 456 1026 462
rect 269 448 318 453
rect -103 440 93 447
rect -104 432 165 437
rect 313 394 318 448
rect 1020 445 1027 452
rect 350 402 355 407
rect 313 388 363 394
rect 1141 366 1221 370
rect 960 362 968 366
rect 268 355 346 360
rect 960 358 1038 362
rect -103 347 81 354
rect 1021 350 1025 354
rect -103 339 165 344
rect 1153 312 1160 314
rect 1153 308 1181 312
rect 1171 302 1181 308
rect 213 297 355 302
rect 1141 266 1215 270
rect 980 258 1038 262
rect 261 254 294 258
rect 289 251 294 254
rect 960 254 968 257
rect 960 250 1031 254
rect 960 249 968 250
rect 257 179 312 183
rect 307 178 312 179
rect 1144 168 1211 172
rect 1001 160 1038 164
rect 1001 158 1007 160
rect 1017 152 1023 157
rect 351 112 357 149
rect 459 116 466 123
rect 277 108 357 112
rect 307 99 362 105
rect 1037 92 1041 121
rect 298 83 393 90
rect 924 89 1041 92
rect 866 82 876 83
rect 866 76 1023 82
rect 866 75 876 76
rect 277 68 367 74
rect 289 57 369 60
rect 289 54 350 57
rect 355 54 369 57
rect 990 45 1000 56
rect 326 33 331 34
rect 282 29 331 33
rect 547 -15 553 19
rect 599 6 605 19
rect 725 10 733 18
rect 936 16 941 29
rect 599 -1 959 6
rect 990 -15 999 45
rect 547 -22 999 -15
<< m2contact >>
rect 363 388 371 394
rect 972 258 980 263
<< metal2 >>
rect 363 -4 371 388
rect 972 -4 980 258
rect 363 -12 980 -4
<< m3contact >>
rect 277 632 283 637
rect 298 540 304 545
rect 326 509 331 514
rect 340 500 345 505
rect 350 402 355 407
rect 340 355 345 360
rect 213 297 218 302
rect 350 297 355 302
rect 289 251 294 258
rect 307 178 312 183
rect 307 99 312 105
rect 298 83 303 90
rect 277 68 283 74
rect 289 54 294 60
rect 326 29 331 34
rect 866 75 876 83
rect 1001 158 1007 164
rect 1017 152 1023 157
rect 1017 76 1023 82
<< metal3 >>
rect -103 297 213 302
rect 277 74 283 632
rect 289 60 294 251
rect 298 90 303 540
rect 307 105 312 178
rect 326 34 331 509
rect 340 361 345 500
rect 340 360 346 361
rect 345 355 346 360
rect 340 46 346 355
rect 350 302 354 402
rect 350 64 355 297
rect 800 75 866 82
rect 800 64 808 75
rect 1001 71 1007 158
rect 1017 82 1023 152
rect 350 57 808 64
rect 815 65 1007 71
rect 815 51 821 65
rect 518 46 821 51
rect 340 45 821 46
rect 340 39 525 45
<< m4contact >>
rect 276 645 283 652
rect 298 606 307 614
rect 1020 456 1026 462
rect 1020 445 1027 452
rect 960 358 968 366
rect 1021 350 1026 355
rect 1153 308 1160 314
rect 725 10 733 18
<< metal4 >>
rect 283 645 1024 652
rect 307 613 411 614
rect 307 606 968 613
rect 382 605 634 606
rect 598 404 605 412
rect 960 366 968 606
rect 1020 462 1024 645
rect 1020 409 1025 445
rect 1020 406 1197 409
rect 1021 312 1025 350
rect 1021 308 1153 312
rect 1190 43 1197 406
rect 1005 35 1197 43
rect 725 -26 733 10
rect 1005 -26 1013 35
rect 725 -33 1013 -26
<< m5contact >>
rect 459 116 466 123
rect 936 16 941 23
rect 232 0 238 7
<< metal5 >>
rect 459 7 465 116
rect 941 16 1219 23
rect 238 0 465 7
<< m6contact >>
rect 938 559 946 567
rect 1171 302 1181 312
rect 960 249 968 257
rect 990 45 1000 56
rect 954 -1 962 8
<< metal6 >>
rect 946 559 1016 567
rect 1005 493 1016 559
rect 954 249 960 257
rect 954 8 963 249
rect 1175 56 1181 302
rect 1000 47 1181 56
rect 962 -1 963 8
use propgen  propgen_0
timestamp 1638739068
transform 1 0 151 0 1 583
box -151 -583 133 87
use cla  cla_0
timestamp 1638764848
transform 1 0 453 0 1 461
box -108 -451 503 136
use sumblock  sumblock_0
timestamp 1638747933
transform 1 0 1023 0 1 415
box -38 -296 124 87
<< labels >>
rlabel metal1 -102 624 119 631 1 a3
rlabel metal1 -103 616 165 621 1 b3
rlabel metal1 -103 524 165 529 1 b2
rlabel metal1 -103 432 165 437 1 b1
rlabel metal1 -103 339 165 344 1 b0
rlabel space -102 532 106 539 1 a2
rlabel metal1 -103 440 93 447 1 a1
rlabel metal1 -103 347 81 354 1 a0
rlabel space -103 296 0 302 1 c_in
rlabel metal1 1203 168 1211 172 1 sum0
rlabel metal1 1202 266 1215 270 1 sum1
rlabel metal1 1208 366 1221 370 1 sum2
rlabel metal1 1207 464 1219 468 1 sum3
rlabel space 1202 15 1220 23 1 carry3
rlabel space 153 662 166 670 5 vdd
rlabel space 160 624 168 628 1 a3
rlabel space 159 616 167 620 1 b3
rlabel metal1 262 632 283 637 1 p3
rlabel space 151 583 166 591 1 gnd
rlabel space 151 570 166 578 1 vdd
rlabel space 153 532 166 536 1 a2
rlabel metal1 154 524 165 529 1 b2
rlabel space 153 491 166 499 1 gnd
rlabel metal1 262 540 277 545 1 p2
rlabel metal1 262 632 276 637 1 p3
rlabel metal1 262 540 304 545 1 p2
rlabel space 152 478 166 486 1 vdd
rlabel space 153 440 165 444 1 a1
rlabel metal1 153 432 165 437 1 b1
rlabel space 153 399 166 407 1 gnd
rlabel space 262 448 276 453 1 p1
rlabel space 152 385 166 393 1 vdd
rlabel space 152 347 160 351 1 a0
rlabel metal1 154 339 165 344 1 b0
rlabel space 262 355 276 360 1 p0
rlabel space 152 306 166 314 1 gnd
rlabel space 149 282 176 291 1 vdd
rlabel space 154 253 170 258 1 a3
rlabel space 155 242 172 249 1 b3
rlabel space 155 225 177 233 1 gnd
rlabel space 156 207 175 216 1 vdd
rlabel space 230 254 248 258 1 g3
rlabel space 158 179 169 184 1 a2
rlabel space 157 167 171 174 1 b2
rlabel space 228 179 255 183 1 g2
rlabel space 157 150 176 158 1 gnd
rlabel space 158 132 175 141 1 vdd
rlabel space 157 104 169 109 1 a1
rlabel space 156 92 171 99 1 b1
rlabel space 156 75 176 83 1 gnd
rlabel space 229 104 256 108 1 g1
rlabel space 158 57 175 66 1 vdd
rlabel space 155 29 169 34 1 a0
rlabel space 154 16 171 24 1 b0
rlabel space 155 0 176 8 1 gnd
rlabel space 229 29 254 33 1 g0
<< end >>
