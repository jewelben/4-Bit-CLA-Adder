* SPICE3 file created from test.ext - technology: scmos

.include TSMC_180nm.txt
.param SUPPLY = 1.8
.option scale=0.09u
.global gnd vdd

VDS vdd gnd 'SUPPLY'
vin1 A gnd pulse 1.8 0 0ns 100ps 100ps 9.9ns 20ns
vin2 B gnd pulse 1.8 0 0ns 100ps 100ps 19.9ns 40ns
vin3 C gnd pulse 1.8 0 0ns 100ps 100ps 39.9ns 80ns
vin4 D gnd pulse 1.8 0 0ns 100ps 100ps 79.9ns 160ns


M1000 VDD 2and_0/B 2and_0/a_13_5# VDD  pfet w=6 l=2
+  ad=252 pd=180 as=48 ps=28
M1001 2or_0/A 2and_0/a_13_5# GND Gnd nfet w=4 l=2
+  ad=20 pd=18 as=140 ps=126
M1002 2and_0/a_13_5# 2and_0/A VDD VDD  pfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1003 2or_0/A 2and_0/a_13_5# VDD VDD  pfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1004 2and_0/a_13_5# 2and_0/B VDD  Gnd nfet w=4 l=2
+  ad=24 pd=20 as=32 ps=24
M1005 VDD  2and_0/A GND Gnd nfet w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1006 VDD 2and_1/B 2and_1/a_13_5# VDD  pfet w=6 l=2
+  ad=0 pd=0 as=48 ps=28
M1007 OUT1 2and_1/a_13_5# GND Gnd nfet w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1008 2and_1/a_13_5# 2and_1/A VDD VDD  pfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1009 OUT1 2and_1/a_13_5# VDD VDD  pfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1010 2and_1/a_13_5# 2and_1/B 2and_1/a_13_n25# Gnd nfet w=4 l=2
+  ad=24 pd=20 as=32 ps=24
M1011 2and_1/a_13_n25# 2and_1/A GND Gnd nfet w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1012 OUTPUT 2or_0/NOR VDD VDD  pfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1013 GND OUT1 2or_0/NOR Gnd nfet w=4 l=2
+  ad=0 pd=0 as=32 ps=24
M1014 2or_0/NOR OUT1 2or_0/a_0_6# VDD  pfet w=6 l=2
+  ad=30 pd=22 as=48 ps=28
M1015 OUTPUT 2or_0/NOR GND Gnd nfet w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1016 2or_0/a_0_6# 2or_0/A VDD VDD  pfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1017 2or_0/NOR 2or_0/A GND Gnd nfet w=4 l=2
+  ad=0 pd=0 as=0 ps=0
C0 2and_1/a_13_5# 2and_1/A 0.04fF
C1 VDD 2or_0/NOR 0.04fF
C2 OUT1 VDD  0.06fF
C3 2and_0/a_13_5# 2and_0/B 0.17fF
C4 2or_0/NOR GND 0.13fF
C5 2and_1/B 2and_1/A 0.24fF
C6 2and_1/a_13_5# VDD  0.08fF
C7 2and_0/a_13_5# VDD  0.08fF
C8 2or_0/A VDD  0.06fF
C9 OUT1 2and_1/a_13_5# 0.05fF
C10 2and_0/a_13_5# 2and_0/A 0.04fF
C11 2and_1/a_13_5# VDD  0.02fF
C12 2and_0/a_13_5# VDD  0.02fF
C13 2and_0/B 2and_0/A 0.26fF
C14 VDD VDD  0.06fF
C15 2or_0/A 2and_0/a_13_5# 0.05fF
C16 2and_1/B VDD  0.08fF
C17 2and_0/B VDD  0.08fF
C18 2or_0/NOR VDD  0.09fF
C19 VDD 2and_1/a_13_5# 0.09fF
C20 2and_1/a_13_5# GND 0.02fF
C21 2and_1/A VDD  0.08fF
C22 2and_0/A VDD  0.08fF
C23 OUT1 VDD  0.03fF
C24 OUTPUT VDD 0.06fF
C25 VDD 2and_0/a_13_5# 0.09fF
C26 2or_0/A VDD  0.03fF
C27 OUTPUT GND 0.06fF
C28 GND 2and_0/a_13_5# 0.02fF
C29 2and_1/B GND 0.03fF
C30 OUTPUT 2or_0/NOR 0.05fF
C31 VDD 2and_0/B 0.03fF
C32 OUT1 2or_0/A 0.43fF
C33 GND 2and_0/B 0.03fF
C34 m5_n1_n2# VDD 0.09fF
C35 VDD VDD  0.03fF
C36 VDD 2and_0/A 0.03fF
C37 m5_n1_n2# GND 0.06fF
C38 VDD VDD  0.03fF
C39 VDD OUT1 0.06fF
C40 VDD VDD  0.06fF
C41 OUT1 GND 0.06fF
C42 VDD VDD  0.06fF
C43 OUTPUT VDD  0.03fF
C44 2or_0/NOR OUT1 0.19fF
C45 VDD 2or_0/A 0.06fF
C46 2or_0/A GND 0.06fF
C47 2and_1/a_13_5# 2and_1/B 0.17fF
C48 m5_n1_n2# Gnd 0.91fF
C49 OUTPUT Gnd 0.22fF
C50 VDD Gnd 1.61fF
C51 2or_0/NOR Gnd 0.35fF
C52 OUT1 Gnd 0.48fF
C53 2or_0/A Gnd 0.35fF
C54 VDD  Gnd 1.03fF
C55 2and_1/a_13_5# Gnd 0.37fF
C56 2and_1/B Gnd 0.34fF
C57 2and_1/A Gnd 0.31fF
C58 VDD  Gnd 0.43fF
C59 VDD  Gnd 0.67fF
C60 GND Gnd 1.14fF
C61 2and_0/a_13_5# Gnd 0.37fF
C62 2and_0/B Gnd 0.34fF
C63 2and_0/A Gnd 0.30fF
C64 VDD  Gnd 0.43fF
C65 VDD  Gnd 0.67fF

.tran 0.05n 160n

.control
run

set color0 = white
set color1 = black

plot v(OUT) v(A)+2 v(B)+4 v(C)+6 v(D)+8


.endc
