magic
tech scmos
timestamp 1638571184
<< metal1 >>
rect -13 61 113 66
rect -13 -12 -9 61
rect 103 51 113 61
rect -3 28 13 32
rect 75 28 91 32
rect -4 19 12 23
rect 87 22 91 28
rect 87 18 101 22
rect 90 11 101 15
rect 153 13 172 17
rect -13 -15 4 -12
rect 90 -44 94 11
rect -2 -48 14 -44
rect 72 -48 94 -44
rect -2 -57 14 -53
rect 154 -71 158 -13
rect 71 -76 160 -71
<< m6contact >>
rect -1 -2 7 6
rect 1 -76 9 -68
<< metal6 >>
rect -10 -2 -1 6
rect -10 -68 -4 -2
rect -10 -76 1 -68
use 2and  2and_0 /media/jewel/SSD/VLSID/Project/Magic/2AND
timestamp 1637099764
transform 1 0 5 0 1 35
box -5 -35 71 29
use 2and  2and_1
timestamp 1637099764
transform 1 0 4 0 1 -41
box -5 -35 71 29
use 2or  2or_0 /media/jewel/SSD/VLSID/Project/Magic/2OR
timestamp 1637169033
transform 1 0 116 0 1 25
box -17 -42 49 29
<< labels >>
rlabel space -3 28 16 32 1 In1
rlabel space -4 19 22 23 1 In2
rlabel space -2 -48 15 -44 1 In3
rlabel space -2 -57 25 -53 1 In4
rlabel metal1 74 -48 94 -44 1 OUT1
rlabel space 72 28 91 32 1 OUT2
rlabel metal1 153 13 172 17 1 OUTPUT
rlabel space -13 61 113 67 5 VDD
rlabel space -10 -76 160 -73 1 GND
<< end >>
